grammar edu:umn:cs:melt:ableJ14:composed:java_sql;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:sql;
imports edu:umn:cs:melt:ableJ14:host only Root_C;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_sql;
} 
