grammar edu:umn:cs:melt:ableJ14:composed:java_complex;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:complex;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_complex;
} 
