grammar edu:umn:cs:melt:ableJ14:composed:java_alone;
exports edu:umn:cs:melt:ableJ14:host;
imports edu:umn:cs:melt:ableJ14:host only Root_C;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_alone;
} 
