grammar edu:umn:cs:melt:ableJ14:composed:java_tables;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:tables;
imports edu:umn:cs:melt:ableJ14:host only Root_C;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_tables;
}
