grammar edu:umn:cs:melt:ableJ14:host;

exports edu:umn:cs:melt:ableJ14:terminals;
exports edu:umn:cs:melt:ableJ14:concretesyntax;
exports edu:umn:cs:melt:ableJ14:abstractsyntax;
exports edu:umn:cs:melt:ableJ14:driver:strict;
exports edu:umn:cs:melt:ableJ14:host:exts:parameterized_expr_block;

import edu:umn:cs:melt:ableJ14:concretesyntax ;

parser hostParse :: Root_C
{
  edu:umn:cs:melt:ableJ14:terminals;
  edu:umn:cs:melt:ableJ14:concretesyntax;
  edu:umn:cs:melt:ableJ14:host:exts:parameterized_expr_block;
}
