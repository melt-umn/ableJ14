grammar edu:umn:cs:melt:ableJ14:composed:java_complex;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:complex;
imports edu:umn:cs:melt:ableJ14:host only Root_C;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_complex;
} 
