grammar edu:umn:cs:melt:ableJ14:composed:java_foreach;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:foreach;
imports edu:umn:cs:melt:ableJ14:host only Root_C;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_foreach;
} 
