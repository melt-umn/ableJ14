grammar edu:umn:cs:melt:ableJ14:composed:java_foreach;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:foreach;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_foreach;
} 
