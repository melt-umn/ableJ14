grammar edu:umn:cs:melt:ableJ14:composed:java_sql;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:sql;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_sql;
} 
