grammar edu:umn:cs:melt:ableJ14:composed:java_pizza;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:pizza:algebraic;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_pizza;
}
