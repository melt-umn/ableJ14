grammar edu:umn:cs:melt:ableJ14:composed:java_autoboxing;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:autoboxing;
parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_autoboxing;
}
