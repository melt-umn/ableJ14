grammar edu:umn:cs:melt:ableJ14:composed:java_rlp;
exports edu:umn:cs:melt:ableJ14:host;
exports edu:umn:cs:melt:ableJ14:exts:rlp;

parser parse :: Root_C {
 edu:umn:cs:melt:ableJ14:composed:java_rlp;
} 
